-----------------------------------------------------------------------
-- Title: Font 5x7
-- Author: zwenergy
-----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity font5x7 is
  port(
    char : in integer range 0 to 37;
    x : in integer range 0 to 4;
    y : in integer range 0 to 6;
    
    clk : in std_logic;
    rst : in std_logic;
    
    charPxl : out std_logic
  );
end entity;

architecture rtl of font5x7 is
type tFontRAM is array( 0 to 37 ) of std_logic_vector( 0 to 34 );
constant font : tFontRAM := 
( "00000000000000000000000000000000000", -- 0, Space
  "01110100011000111111100011000110001", -- 1, A
  "11110100011000111110100011000111110", -- 2, B
  "11111100001000010000100001000011111", -- 3, C
  "11110100011000110001100011000111110", -- 4, D
  "11111100001000011110100001000011111", -- 5, E
  "11111100001000011110100001000010000", -- 6, F
  "01111100001000010011100011000101110", -- 7, G
  "10001100011000111111100011000110001", -- 8, H
  "01110001000010000100001000010001110", -- 9, I
  "11111000010000100001000011000101110", -- 10, J
  "10001100011001011100100101000110001", -- 11, K
  "10000100001000010000100001000011111", -- 12, L
  "10001110111010110001100011000110001", -- 13, M
  "10001110011100110101100111001110001", -- 14, N
  "01110100011000110001100011000101110", -- 15, O
  "11110100011000111110100001000010000", -- 16, P
  "01110100011000101111000010000100001", -- 17, Q
  "11110100011000111110100011000110001", -- 18, R
  "01111100001000001110000010000111110", -- 19, S
  "11111001000010000100001000010000100", -- 20, T
  "10001100011000110001100011000101110", -- 21, U
  "10001100011000101010010100010000100", -- 22, V
  "10001100011000110001100011010101010", -- 23, W
  "10001100010101000100010101000110001", -- 24, X
  "10001100010101000100001000010000100", -- 25, Y
  "11111000010001000100010001000011111", -- 26, Z
  "00100011000010000100001000010001110", -- 27, 1
  "01110100010000100010001000100011111", -- 28, 2
  "01110100010000100110000011000101110", -- 29, 3
  "10000100001010011111001000010000100", -- 30, 4
  "11111100001000001110000010000111110", -- 31, 5
  "01111110001000010110110011000101110", -- 32, 6
  "11111000010001000100010001000010000", -- 33, 7
  "01110100011000101110100011000101110", -- 34, 8
  "01110100011000101111000010000100001", -- 35, 9
  "00000000000000000000000000000000100", -- 36, .
  "00000010000010000010001000100000000"  -- 37, >
  );
begin

  process( clk )  is
  variable offset : integer range 0 to 30;
  variable ind : integer range 0 to 34;
  begin
    if ( rising_edge( clk ) )  then
      if ( rst = '1' ) then
        charPxl <= '0';
      else
        offset := 0;
        case y is
          when 0 => offset := 0;
          when 1 => offset := 5;
          when 2 => offset := 10;
          when 3 => offset := 15;
          when 4 => offset := 20;
          when 5 => offset := 25;
          when 6 => offset := 30;
        end case;
        
        ind := offset + x;
        
        charPxl <= font( char )( ind );
      end if;
    end if;
  
  end process;

end rtl;
